`ifndef add16
  `include "src/add16.v"
`endif

module add16_test;
  reg [15:0] a, b;
  wire [15:0] out;

  add16 u (a, b, out);

  initial begin
    a = 16'b0000000000000000;
    b = 16'b0000000000000000;
    #1;
    assert((a + b) == out);

    a = 16'b0000000000000001;
    b = 16'b0000000000000001;
    #1;
    assert((a + b) == out);

    a = 16'b0000000000000001;
    b = 16'b0000000000000010;
    #1;
    assert((a + b) == out);

    a = 16'b1000000000000001;
    b = 16'b1000000000000001;
    #1;
    assert((a + b) == out);

    a = 16'b1010101010101010;
    b = 16'b0101010101010101;
    #1;
    assert((a + b) == out);

    a = 16'b1111111111111111;
    b = 16'b0000000000000000;
    #1;
    assert((a + b) == out);

    a = 16'b1111111111111111;
    b = 16'b1111111111111111;
    #1;
    assert((a + b) == out);

    a = 16'b1111111100000000;
    b = 16'b0000000011111111;
    #1;
    assert((a + b) == out);

    a = 16'b0010101010010100;
    b = 16'b1010010010010101;
    #1;
    assert((a + b) == out);

    a = 16'b0111111111111111;
    b = 16'b0000000000000001;
    #1;
    assert((a + b) == out);
  end
endmodule;
